

module pipeline_tb ();




endmodule